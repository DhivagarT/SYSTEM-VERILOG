# KERNEL: a=4 b=6 y=10
