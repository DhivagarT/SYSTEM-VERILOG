module sum(add.dut intf);
  
  assign intf.y=intf.a + intf.b;

endmodule
