interface xor_int;
  logic a;
  logic b;
  logic y;
endinterface
