module xor_des(xor_int intrf);
  
  assign intrf.y=intrf.a ^ intrf.b;
  
endmodule
