a=0 b=x y=x
a=0 b=1 y=1
a=1 b=1 y=0
a=1 b=0 y=1
a=1 b=1 y=0
